LIBRARY ieee;
USE ieee.STD_LOGIC_1164.ALL;
USE ieee.NUMERIC_STD.ALL;

PACKAGE ya_uart_pkg IS
  
  CONSTANT C_CLK_FREQ_HZ        : INTEGER := 125000000;
  
  -- Baudrate constants
  CONSTANT C_BAUD_9600_HZ       : INTEGER := 9600;
  CONSTANT C_BAUD_19200_HZ      : INTEGER := 19200;
  CONSTANT C_BAUD_CNT_MAX       : INTEGER := 65535; 
  CONSTANT C_INCREMENT          : INTEGER := 1;

  CONSTANT C_DIV_9600_CYC       : INTEGER := C_CLK_FREQ_HZ / C_BAUD_9600_HZ;
  CONSTANT C_DIV_19200_CYC      : INTEGER := C_CLK_FREQ_HZ / C_BAUD_19200_HZ;

  CONSTANT C_DIV_9600_FULL_MAX  : INTEGER := C_DIV_9600_CYC - 1;
  CONSTANT C_DIV_19200_FULL_MAX : INTEGER := C_DIV_19200_CYC - 1;

  CONSTANT C_DIV_9600_HALF_MAX  : INTEGER := (C_DIV_9600_CYC / 2) - 1;
  CONSTANT C_DIV_19200_HALF_MAX : INTEGER := (C_DIV_19200_CYC / 2) - 1;

  -- Baudrate Testbench  constants
  CONSTANT C_TB_CLK_PERIOD_NS : TIME := 8 ns;
  CONSTANT C_TB_RESET_TIME_NS : TIME := 100 ns;
  CONSTANT C_TB_RUN_TIME_MS   : TIME := 5 ms;

END PACKAGE ya_uart_pkg;