ARCHITECTURE ha_a OF ha_e IS 
BEGIN 

  s_o <= a_i XOR b_i;
  c_o <= a_i AND b_i;
  
END ha_a;
