LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.all;
    USE IEEE.NUMERIC_STD.all;
    
    
ENTITY ha_e IS 
PORT(
  a_i : IN  std_logic;
  b_i : IN  std_logic;
  s_o : OUT std_logic;
  c_o : OUT std_logic
  );
END ha_e;

